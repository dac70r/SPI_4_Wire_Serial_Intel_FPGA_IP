// spi_platform_designer.v

// Generated using ACDS version 23.1 993

`timescale 1 ps / 1 ps
module spi_platform_designer (
		input  wire  clk_clk,                  //               clk.clk
		input  wire  esc_eepdone_input_export, // esc_eepdone_input.export
		input  wire  esc_spi_MISO,             //           esc_spi.MISO
		output wire  esc_spi_MOSI,             //                  .MOSI
		output wire  esc_spi_SCLK,             //                  .SCLK
		output wire  esc_spi_SS_n,             //                  .SS_n
		output wire  esc_spi_cs_export,        //        esc_spi_cs.export
		output wire  led_export,               //               led.export
		input  wire  reset_reset_n             //             reset.reset_n
	);

	wire  [31:0] nios_data_master_readdata;                             // mm_interconnect_0:NIOS_data_master_readdata -> NIOS:d_readdata
	wire         nios_data_master_waitrequest;                          // mm_interconnect_0:NIOS_data_master_waitrequest -> NIOS:d_waitrequest
	wire         nios_data_master_debugaccess;                          // NIOS:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOS_data_master_debugaccess
	wire  [17:0] nios_data_master_address;                              // NIOS:d_address -> mm_interconnect_0:NIOS_data_master_address
	wire   [3:0] nios_data_master_byteenable;                           // NIOS:d_byteenable -> mm_interconnect_0:NIOS_data_master_byteenable
	wire         nios_data_master_read;                                 // NIOS:d_read -> mm_interconnect_0:NIOS_data_master_read
	wire         nios_data_master_write;                                // NIOS:d_write -> mm_interconnect_0:NIOS_data_master_write
	wire  [31:0] nios_data_master_writedata;                            // NIOS:d_writedata -> mm_interconnect_0:NIOS_data_master_writedata
	wire  [31:0] nios_instruction_master_readdata;                      // mm_interconnect_0:NIOS_instruction_master_readdata -> NIOS:i_readdata
	wire         nios_instruction_master_waitrequest;                   // mm_interconnect_0:NIOS_instruction_master_waitrequest -> NIOS:i_waitrequest
	wire  [17:0] nios_instruction_master_address;                       // NIOS:i_address -> mm_interconnect_0:NIOS_instruction_master_address
	wire         nios_instruction_master_read;                          // NIOS:i_read -> mm_interconnect_0:NIOS_instruction_master_read
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_readdata;       // NIOS:debug_mem_slave_readdata -> mm_interconnect_0:NIOS_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios_debug_mem_slave_waitrequest;    // NIOS:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOS_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios_debug_mem_slave_debugaccess;    // mm_interconnect_0:NIOS_debug_mem_slave_debugaccess -> NIOS:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios_debug_mem_slave_address;        // mm_interconnect_0:NIOS_debug_mem_slave_address -> NIOS:debug_mem_slave_address
	wire         mm_interconnect_0_nios_debug_mem_slave_read;           // mm_interconnect_0:NIOS_debug_mem_slave_read -> NIOS:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios_debug_mem_slave_byteenable;     // mm_interconnect_0:NIOS_debug_mem_slave_byteenable -> NIOS:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios_debug_mem_slave_write;          // mm_interconnect_0:NIOS_debug_mem_slave_write -> NIOS:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_writedata;      // mm_interconnect_0:NIOS_debug_mem_slave_writedata -> NIOS:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                   // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                     // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire  [13:0] mm_interconnect_0_ram_s1_address;                      // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                   // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                        // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                    // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                        // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire         mm_interconnect_0_esc_spi_cs_s1_chipselect;            // mm_interconnect_0:ESC_SPI_CS_s1_chipselect -> ESC_SPI_CS:chipselect
	wire  [31:0] mm_interconnect_0_esc_spi_cs_s1_readdata;              // ESC_SPI_CS:readdata -> mm_interconnect_0:ESC_SPI_CS_s1_readdata
	wire   [1:0] mm_interconnect_0_esc_spi_cs_s1_address;               // mm_interconnect_0:ESC_SPI_CS_s1_address -> ESC_SPI_CS:address
	wire         mm_interconnect_0_esc_spi_cs_s1_write;                 // mm_interconnect_0:ESC_SPI_CS_s1_write -> ESC_SPI_CS:write_n
	wire  [31:0] mm_interconnect_0_esc_spi_cs_s1_writedata;             // mm_interconnect_0:ESC_SPI_CS_s1_writedata -> ESC_SPI_CS:writedata
	wire  [31:0] mm_interconnect_0_esc_eepdone_input_s1_readdata;       // ESC_EEPDONE_INPUT:readdata -> mm_interconnect_0:ESC_EEPDONE_INPUT_s1_readdata
	wire   [1:0] mm_interconnect_0_esc_eepdone_input_s1_address;        // mm_interconnect_0:ESC_EEPDONE_INPUT_s1_address -> ESC_EEPDONE_INPUT:address
	wire         mm_interconnect_0_led_s1_chipselect;                   // mm_interconnect_0:LED_s1_chipselect -> LED:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                     // LED:readdata -> mm_interconnect_0:LED_s1_readdata
	wire   [1:0] mm_interconnect_0_led_s1_address;                      // mm_interconnect_0:LED_s1_address -> LED:address
	wire         mm_interconnect_0_led_s1_write;                        // mm_interconnect_0:LED_s1_write -> LED:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                    // mm_interconnect_0:LED_s1_writedata -> LED:writedata
	wire         mm_interconnect_0_esc_spi_spi_control_port_chipselect; // mm_interconnect_0:ESC_SPI_spi_control_port_chipselect -> ESC_SPI:spi_select
	wire  [15:0] mm_interconnect_0_esc_spi_spi_control_port_readdata;   // ESC_SPI:data_to_cpu -> mm_interconnect_0:ESC_SPI_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_esc_spi_spi_control_port_address;    // mm_interconnect_0:ESC_SPI_spi_control_port_address -> ESC_SPI:mem_addr
	wire         mm_interconnect_0_esc_spi_spi_control_port_read;       // mm_interconnect_0:ESC_SPI_spi_control_port_read -> ESC_SPI:read_n
	wire         mm_interconnect_0_esc_spi_spi_control_port_write;      // mm_interconnect_0:ESC_SPI_spi_control_port_write -> ESC_SPI:write_n
	wire  [15:0] mm_interconnect_0_esc_spi_spi_control_port_writedata;  // mm_interconnect_0:ESC_SPI_spi_control_port_writedata -> ESC_SPI:data_from_cpu
	wire         irq_mapper_receiver0_irq;                              // ESC_SPI:irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios_irq_irq;                                          // irq_mapper:sender_irq -> NIOS:irq
	wire         rst_controller_reset_out_reset;                        // rst_controller:reset_out -> [ESC_EEPDONE_INPUT:reset_n, ESC_SPI:reset_n, ESC_SPI_CS:reset_n, LED:reset_n, NIOS:reset_n, RAM:reset, irq_mapper:reset, mm_interconnect_0:NIOS_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                    // rst_controller:reset_req -> [NIOS:reset_req, RAM:reset_req, rst_translator:reset_req_in]

	spi_platform_designer_ESC_EEPDONE_INPUT esc_eepdone_input (
		.clk      (clk_clk),                                         //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address  (mm_interconnect_0_esc_eepdone_input_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_esc_eepdone_input_s1_readdata), //                    .readdata
		.in_port  (esc_eepdone_input_export)                         // external_connection.export
	);

	spi_platform_designer_ESC_SPI esc_spi (
		.clk           (clk_clk),                                               //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                       //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_esc_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_esc_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_esc_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_esc_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_esc_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_esc_spi_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver0_irq),                              //              irq.irq
		.MISO          (esc_spi_MISO),                                          //         external.export
		.MOSI          (esc_spi_MOSI),                                          //                 .export
		.SCLK          (esc_spi_SCLK),                                          //                 .export
		.SS_n          (esc_spi_SS_n)                                           //                 .export
	);

	spi_platform_designer_ESC_SPI_CS esc_spi_cs (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_esc_spi_cs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_esc_spi_cs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_esc_spi_cs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_esc_spi_cs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_esc_spi_cs_s1_readdata),   //                    .readdata
		.out_port   (esc_spi_cs_export)                           // external_connection.export
	);

	spi_platform_designer_LED led (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_export)                           // external_connection.export
	);

	spi_platform_designer_NIOS nios (
		.clk                                 (clk_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                    //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                 //                          .reset_req
		.d_address                           (nios_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_data_master_read),                              //                          .read
		.d_readdata                          (nios_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_data_master_write),                             //                          .write
		.d_writedata                         (nios_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                   //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                    // custom_instruction_master.readra
	);

	spi_platform_designer_RAM ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	spi_platform_designer_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                          (clk_clk),                                               //                        clk_0_clk.clk
		.NIOS_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                        // NIOS_reset_reset_bridge_in_reset.reset
		.NIOS_data_master_address               (nios_data_master_address),                              //                 NIOS_data_master.address
		.NIOS_data_master_waitrequest           (nios_data_master_waitrequest),                          //                                 .waitrequest
		.NIOS_data_master_byteenable            (nios_data_master_byteenable),                           //                                 .byteenable
		.NIOS_data_master_read                  (nios_data_master_read),                                 //                                 .read
		.NIOS_data_master_readdata              (nios_data_master_readdata),                             //                                 .readdata
		.NIOS_data_master_write                 (nios_data_master_write),                                //                                 .write
		.NIOS_data_master_writedata             (nios_data_master_writedata),                            //                                 .writedata
		.NIOS_data_master_debugaccess           (nios_data_master_debugaccess),                          //                                 .debugaccess
		.NIOS_instruction_master_address        (nios_instruction_master_address),                       //          NIOS_instruction_master.address
		.NIOS_instruction_master_waitrequest    (nios_instruction_master_waitrequest),                   //                                 .waitrequest
		.NIOS_instruction_master_read           (nios_instruction_master_read),                          //                                 .read
		.NIOS_instruction_master_readdata       (nios_instruction_master_readdata),                      //                                 .readdata
		.ESC_EEPDONE_INPUT_s1_address           (mm_interconnect_0_esc_eepdone_input_s1_address),        //             ESC_EEPDONE_INPUT_s1.address
		.ESC_EEPDONE_INPUT_s1_readdata          (mm_interconnect_0_esc_eepdone_input_s1_readdata),       //                                 .readdata
		.ESC_SPI_spi_control_port_address       (mm_interconnect_0_esc_spi_spi_control_port_address),    //         ESC_SPI_spi_control_port.address
		.ESC_SPI_spi_control_port_write         (mm_interconnect_0_esc_spi_spi_control_port_write),      //                                 .write
		.ESC_SPI_spi_control_port_read          (mm_interconnect_0_esc_spi_spi_control_port_read),       //                                 .read
		.ESC_SPI_spi_control_port_readdata      (mm_interconnect_0_esc_spi_spi_control_port_readdata),   //                                 .readdata
		.ESC_SPI_spi_control_port_writedata     (mm_interconnect_0_esc_spi_spi_control_port_writedata),  //                                 .writedata
		.ESC_SPI_spi_control_port_chipselect    (mm_interconnect_0_esc_spi_spi_control_port_chipselect), //                                 .chipselect
		.ESC_SPI_CS_s1_address                  (mm_interconnect_0_esc_spi_cs_s1_address),               //                    ESC_SPI_CS_s1.address
		.ESC_SPI_CS_s1_write                    (mm_interconnect_0_esc_spi_cs_s1_write),                 //                                 .write
		.ESC_SPI_CS_s1_readdata                 (mm_interconnect_0_esc_spi_cs_s1_readdata),              //                                 .readdata
		.ESC_SPI_CS_s1_writedata                (mm_interconnect_0_esc_spi_cs_s1_writedata),             //                                 .writedata
		.ESC_SPI_CS_s1_chipselect               (mm_interconnect_0_esc_spi_cs_s1_chipselect),            //                                 .chipselect
		.LED_s1_address                         (mm_interconnect_0_led_s1_address),                      //                           LED_s1.address
		.LED_s1_write                           (mm_interconnect_0_led_s1_write),                        //                                 .write
		.LED_s1_readdata                        (mm_interconnect_0_led_s1_readdata),                     //                                 .readdata
		.LED_s1_writedata                       (mm_interconnect_0_led_s1_writedata),                    //                                 .writedata
		.LED_s1_chipselect                      (mm_interconnect_0_led_s1_chipselect),                   //                                 .chipselect
		.NIOS_debug_mem_slave_address           (mm_interconnect_0_nios_debug_mem_slave_address),        //             NIOS_debug_mem_slave.address
		.NIOS_debug_mem_slave_write             (mm_interconnect_0_nios_debug_mem_slave_write),          //                                 .write
		.NIOS_debug_mem_slave_read              (mm_interconnect_0_nios_debug_mem_slave_read),           //                                 .read
		.NIOS_debug_mem_slave_readdata          (mm_interconnect_0_nios_debug_mem_slave_readdata),       //                                 .readdata
		.NIOS_debug_mem_slave_writedata         (mm_interconnect_0_nios_debug_mem_slave_writedata),      //                                 .writedata
		.NIOS_debug_mem_slave_byteenable        (mm_interconnect_0_nios_debug_mem_slave_byteenable),     //                                 .byteenable
		.NIOS_debug_mem_slave_waitrequest       (mm_interconnect_0_nios_debug_mem_slave_waitrequest),    //                                 .waitrequest
		.NIOS_debug_mem_slave_debugaccess       (mm_interconnect_0_nios_debug_mem_slave_debugaccess),    //                                 .debugaccess
		.RAM_s1_address                         (mm_interconnect_0_ram_s1_address),                      //                           RAM_s1.address
		.RAM_s1_write                           (mm_interconnect_0_ram_s1_write),                        //                                 .write
		.RAM_s1_readdata                        (mm_interconnect_0_ram_s1_readdata),                     //                                 .readdata
		.RAM_s1_writedata                       (mm_interconnect_0_ram_s1_writedata),                    //                                 .writedata
		.RAM_s1_byteenable                      (mm_interconnect_0_ram_s1_byteenable),                   //                                 .byteenable
		.RAM_s1_chipselect                      (mm_interconnect_0_ram_s1_chipselect),                   //                                 .chipselect
		.RAM_s1_clken                           (mm_interconnect_0_ram_s1_clken)                         //                                 .clken
	);

	spi_platform_designer_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios_irq_irq)                    //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
