// spi_platform_designer.v

// Generated using ACDS version 23.1 991

`timescale 1 ps / 1 ps
module spi_platform_designer (
		input  wire  clk_clk,              //           clk.clk
		input  wire  reset_reset_n,        //         reset.reset_n
		input  wire  spi_pin_MISO,         //       spi_pin.MISO
		output wire  spi_pin_MOSI,         //              .MOSI
		output wire  spi_pin_SCLK,         //              .SCLK
		output wire  spi_pin_SS_n,         //              .SS_n
		output wire  spi_ss_manual_export  // spi_ss_manual.export
	);

	wire  [31:0] nios_data_master_readdata;                             // mm_interconnect_0:NIOS_data_master_readdata -> NIOS:d_readdata
	wire         nios_data_master_waitrequest;                          // mm_interconnect_0:NIOS_data_master_waitrequest -> NIOS:d_waitrequest
	wire         nios_data_master_debugaccess;                          // NIOS:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOS_data_master_debugaccess
	wire  [17:0] nios_data_master_address;                              // NIOS:d_address -> mm_interconnect_0:NIOS_data_master_address
	wire   [3:0] nios_data_master_byteenable;                           // NIOS:d_byteenable -> mm_interconnect_0:NIOS_data_master_byteenable
	wire         nios_data_master_read;                                 // NIOS:d_read -> mm_interconnect_0:NIOS_data_master_read
	wire         nios_data_master_write;                                // NIOS:d_write -> mm_interconnect_0:NIOS_data_master_write
	wire  [31:0] nios_data_master_writedata;                            // NIOS:d_writedata -> mm_interconnect_0:NIOS_data_master_writedata
	wire  [31:0] nios_instruction_master_readdata;                      // mm_interconnect_0:NIOS_instruction_master_readdata -> NIOS:i_readdata
	wire         nios_instruction_master_waitrequest;                   // mm_interconnect_0:NIOS_instruction_master_waitrequest -> NIOS:i_waitrequest
	wire  [17:0] nios_instruction_master_address;                       // NIOS:i_address -> mm_interconnect_0:NIOS_instruction_master_address
	wire         nios_instruction_master_read;                          // NIOS:i_read -> mm_interconnect_0:NIOS_instruction_master_read
	wire         mm_interconnect_0_debug_avalon_jtag_slave_chipselect;  // mm_interconnect_0:DEBUG_avalon_jtag_slave_chipselect -> DEBUG:av_chipselect
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_readdata;    // DEBUG:av_readdata -> mm_interconnect_0:DEBUG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_debug_avalon_jtag_slave_waitrequest; // DEBUG:av_waitrequest -> mm_interconnect_0:DEBUG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_debug_avalon_jtag_slave_address;     // mm_interconnect_0:DEBUG_avalon_jtag_slave_address -> DEBUG:av_address
	wire         mm_interconnect_0_debug_avalon_jtag_slave_read;        // mm_interconnect_0:DEBUG_avalon_jtag_slave_read -> DEBUG:av_read_n
	wire         mm_interconnect_0_debug_avalon_jtag_slave_write;       // mm_interconnect_0:DEBUG_avalon_jtag_slave_write -> DEBUG:av_write_n
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_writedata;   // mm_interconnect_0:DEBUG_avalon_jtag_slave_writedata -> DEBUG:av_writedata
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_readdata;       // NIOS:debug_mem_slave_readdata -> mm_interconnect_0:NIOS_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios_debug_mem_slave_waitrequest;    // NIOS:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOS_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios_debug_mem_slave_debugaccess;    // mm_interconnect_0:NIOS_debug_mem_slave_debugaccess -> NIOS:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios_debug_mem_slave_address;        // mm_interconnect_0:NIOS_debug_mem_slave_address -> NIOS:debug_mem_slave_address
	wire         mm_interconnect_0_nios_debug_mem_slave_read;           // mm_interconnect_0:NIOS_debug_mem_slave_read -> NIOS:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios_debug_mem_slave_byteenable;     // mm_interconnect_0:NIOS_debug_mem_slave_byteenable -> NIOS:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios_debug_mem_slave_write;          // mm_interconnect_0:NIOS_debug_mem_slave_write -> NIOS:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_writedata;      // mm_interconnect_0:NIOS_debug_mem_slave_writedata -> NIOS:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                   // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                     // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire  [13:0] mm_interconnect_0_ram_s1_address;                      // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                   // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                        // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                    // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                        // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire         mm_interconnect_0_spi_ss_manual_s1_chipselect;         // mm_interconnect_0:SPI_SS_MANUAL_s1_chipselect -> SPI_SS_MANUAL:chipselect
	wire  [31:0] mm_interconnect_0_spi_ss_manual_s1_readdata;           // SPI_SS_MANUAL:readdata -> mm_interconnect_0:SPI_SS_MANUAL_s1_readdata
	wire   [1:0] mm_interconnect_0_spi_ss_manual_s1_address;            // mm_interconnect_0:SPI_SS_MANUAL_s1_address -> SPI_SS_MANUAL:address
	wire         mm_interconnect_0_spi_ss_manual_s1_write;              // mm_interconnect_0:SPI_SS_MANUAL_s1_write -> SPI_SS_MANUAL:write_n
	wire  [31:0] mm_interconnect_0_spi_ss_manual_s1_writedata;          // mm_interconnect_0:SPI_SS_MANUAL_s1_writedata -> SPI_SS_MANUAL:writedata
	wire         mm_interconnect_0_spi_spi_control_port_chipselect;     // mm_interconnect_0:SPI_spi_control_port_chipselect -> SPI:spi_select
	wire  [15:0] mm_interconnect_0_spi_spi_control_port_readdata;       // SPI:data_to_cpu -> mm_interconnect_0:SPI_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_spi_control_port_address;        // mm_interconnect_0:SPI_spi_control_port_address -> SPI:mem_addr
	wire         mm_interconnect_0_spi_spi_control_port_read;           // mm_interconnect_0:SPI_spi_control_port_read -> SPI:read_n
	wire         mm_interconnect_0_spi_spi_control_port_write;          // mm_interconnect_0:SPI_spi_control_port_write -> SPI:write_n
	wire  [15:0] mm_interconnect_0_spi_spi_control_port_writedata;      // mm_interconnect_0:SPI_spi_control_port_writedata -> SPI:data_from_cpu
	wire         irq_mapper_receiver0_irq;                              // SPI:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                              // DEBUG:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios_irq_irq;                                          // irq_mapper:sender_irq -> NIOS:irq
	wire         rst_controller_reset_out_reset;                        // rst_controller:reset_out -> [DEBUG:rst_n, NIOS:reset_n, RAM:reset, SPI:reset_n, SPI_SS_MANUAL:reset_n, irq_mapper:reset, mm_interconnect_0:NIOS_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                    // rst_controller:reset_req -> [NIOS:reset_req, RAM:reset_req, rst_translator:reset_req_in]

	spi_platform_designer_DEBUG debug (
		.clk            (clk_clk),                                               //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_debug_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_debug_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_debug_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_debug_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_debug_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                               //               irq.irq
	);

	spi_platform_designer_NIOS nios (
		.clk                                 (clk_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                    //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                 //                          .reset_req
		.d_address                           (nios_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_data_master_read),                              //                          .read
		.d_readdata                          (nios_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_data_master_write),                             //                          .write
		.d_writedata                         (nios_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                   //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                    // custom_instruction_master.readra
	);

	spi_platform_designer_RAM ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	spi_platform_designer_SPI spi (
		.clk           (clk_clk),                                           //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                   //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver0_irq),                          //              irq.irq
		.MISO          (spi_pin_MISO),                                      //         external.export
		.MOSI          (spi_pin_MOSI),                                      //                 .export
		.SCLK          (spi_pin_SCLK),                                      //                 .export
		.SS_n          (spi_pin_SS_n)                                       //                 .export
	);

	spi_platform_designer_SPI_SS_MANUAL spi_ss_manual (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_spi_ss_manual_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_spi_ss_manual_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_spi_ss_manual_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_spi_ss_manual_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_spi_ss_manual_s1_readdata),   //                    .readdata
		.out_port   (spi_ss_manual_export)                           // external_connection.export
	);

	spi_platform_designer_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                          (clk_clk),                                               //                        clk_0_clk.clk
		.NIOS_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                        // NIOS_reset_reset_bridge_in_reset.reset
		.NIOS_data_master_address               (nios_data_master_address),                              //                 NIOS_data_master.address
		.NIOS_data_master_waitrequest           (nios_data_master_waitrequest),                          //                                 .waitrequest
		.NIOS_data_master_byteenable            (nios_data_master_byteenable),                           //                                 .byteenable
		.NIOS_data_master_read                  (nios_data_master_read),                                 //                                 .read
		.NIOS_data_master_readdata              (nios_data_master_readdata),                             //                                 .readdata
		.NIOS_data_master_write                 (nios_data_master_write),                                //                                 .write
		.NIOS_data_master_writedata             (nios_data_master_writedata),                            //                                 .writedata
		.NIOS_data_master_debugaccess           (nios_data_master_debugaccess),                          //                                 .debugaccess
		.NIOS_instruction_master_address        (nios_instruction_master_address),                       //          NIOS_instruction_master.address
		.NIOS_instruction_master_waitrequest    (nios_instruction_master_waitrequest),                   //                                 .waitrequest
		.NIOS_instruction_master_read           (nios_instruction_master_read),                          //                                 .read
		.NIOS_instruction_master_readdata       (nios_instruction_master_readdata),                      //                                 .readdata
		.DEBUG_avalon_jtag_slave_address        (mm_interconnect_0_debug_avalon_jtag_slave_address),     //          DEBUG_avalon_jtag_slave.address
		.DEBUG_avalon_jtag_slave_write          (mm_interconnect_0_debug_avalon_jtag_slave_write),       //                                 .write
		.DEBUG_avalon_jtag_slave_read           (mm_interconnect_0_debug_avalon_jtag_slave_read),        //                                 .read
		.DEBUG_avalon_jtag_slave_readdata       (mm_interconnect_0_debug_avalon_jtag_slave_readdata),    //                                 .readdata
		.DEBUG_avalon_jtag_slave_writedata      (mm_interconnect_0_debug_avalon_jtag_slave_writedata),   //                                 .writedata
		.DEBUG_avalon_jtag_slave_waitrequest    (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest), //                                 .waitrequest
		.DEBUG_avalon_jtag_slave_chipselect     (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),  //                                 .chipselect
		.NIOS_debug_mem_slave_address           (mm_interconnect_0_nios_debug_mem_slave_address),        //             NIOS_debug_mem_slave.address
		.NIOS_debug_mem_slave_write             (mm_interconnect_0_nios_debug_mem_slave_write),          //                                 .write
		.NIOS_debug_mem_slave_read              (mm_interconnect_0_nios_debug_mem_slave_read),           //                                 .read
		.NIOS_debug_mem_slave_readdata          (mm_interconnect_0_nios_debug_mem_slave_readdata),       //                                 .readdata
		.NIOS_debug_mem_slave_writedata         (mm_interconnect_0_nios_debug_mem_slave_writedata),      //                                 .writedata
		.NIOS_debug_mem_slave_byteenable        (mm_interconnect_0_nios_debug_mem_slave_byteenable),     //                                 .byteenable
		.NIOS_debug_mem_slave_waitrequest       (mm_interconnect_0_nios_debug_mem_slave_waitrequest),    //                                 .waitrequest
		.NIOS_debug_mem_slave_debugaccess       (mm_interconnect_0_nios_debug_mem_slave_debugaccess),    //                                 .debugaccess
		.RAM_s1_address                         (mm_interconnect_0_ram_s1_address),                      //                           RAM_s1.address
		.RAM_s1_write                           (mm_interconnect_0_ram_s1_write),                        //                                 .write
		.RAM_s1_readdata                        (mm_interconnect_0_ram_s1_readdata),                     //                                 .readdata
		.RAM_s1_writedata                       (mm_interconnect_0_ram_s1_writedata),                    //                                 .writedata
		.RAM_s1_byteenable                      (mm_interconnect_0_ram_s1_byteenable),                   //                                 .byteenable
		.RAM_s1_chipselect                      (mm_interconnect_0_ram_s1_chipselect),                   //                                 .chipselect
		.RAM_s1_clken                           (mm_interconnect_0_ram_s1_clken),                        //                                 .clken
		.SPI_spi_control_port_address           (mm_interconnect_0_spi_spi_control_port_address),        //             SPI_spi_control_port.address
		.SPI_spi_control_port_write             (mm_interconnect_0_spi_spi_control_port_write),          //                                 .write
		.SPI_spi_control_port_read              (mm_interconnect_0_spi_spi_control_port_read),           //                                 .read
		.SPI_spi_control_port_readdata          (mm_interconnect_0_spi_spi_control_port_readdata),       //                                 .readdata
		.SPI_spi_control_port_writedata         (mm_interconnect_0_spi_spi_control_port_writedata),      //                                 .writedata
		.SPI_spi_control_port_chipselect        (mm_interconnect_0_spi_spi_control_port_chipselect),     //                                 .chipselect
		.SPI_SS_MANUAL_s1_address               (mm_interconnect_0_spi_ss_manual_s1_address),            //                 SPI_SS_MANUAL_s1.address
		.SPI_SS_MANUAL_s1_write                 (mm_interconnect_0_spi_ss_manual_s1_write),              //                                 .write
		.SPI_SS_MANUAL_s1_readdata              (mm_interconnect_0_spi_ss_manual_s1_readdata),           //                                 .readdata
		.SPI_SS_MANUAL_s1_writedata             (mm_interconnect_0_spi_ss_manual_s1_writedata),          //                                 .writedata
		.SPI_SS_MANUAL_s1_chipselect            (mm_interconnect_0_spi_ss_manual_s1_chipselect)          //                                 .chipselect
	);

	spi_platform_designer_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios_irq_irq)                    //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
